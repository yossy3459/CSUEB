`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/24/2017 11:12:22 AM
// Design Name: 
// Module Name: shape
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module shape(
    input [4:0] clockCount,
    input [3:0] shapeCount,
    input [8:0] x,
    output [7:0] DB
    );
endmodule
