`timescale 1ns / 1ps
module topmodule(
    input Clk,
    input Rst,
    input [1:0] Fsel,
    input [2:0] Fr,
    output [7:0] DB,
    output CS,
    output WR,
    output AB,
    output PD,
    output LDAC,
    output CLR,
    output VDD,
    output REFIN,
    output VoutA,
    output VoutB,
    output DGND
    );
    
    
    
endmodule