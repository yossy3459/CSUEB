`timescale 1ns / 1ps

module dataCreator(
    input Rst,
    input [1:0] Fsel,
    input dbClock,
    output [7:0] DB
    );
    
    reg [7:0] DB;
    reg [8:0] horizontalCount;
    reg upDownFlag;        // 0 => up, 1 => down
    reg squareInitFlag;

    
    always @( negedge dbClock or negedge Rst ) begin
        if (!Rst) begin
            DB <= 0;
            upDownFlag <= 0;
            horizontalCount <= 0;
        end
        else begin
        case ( Fsel ) 
            // sin
            2'b00: 
                begin 
                    case ( horizontalCount ) 
                    0	 : DB <=	127	   ;
                    1    : DB <=    129    ;
                    2    : DB <=    130    ;
                    3    : DB <=    132    ;
                    4    : DB <=    133    ;
                    5    : DB <=    135    ;
                    6    : DB <=    136    ;
                    7    : DB <=    138    ;
                    8    : DB <=    140    ;
                    9    : DB <=    141    ;
                    10    : DB <=    143    ;
                    11    : DB <=    144    ;
                    12    : DB <=    146    ;
                    13    : DB <=    147    ;
                    14    : DB <=    149    ;
                    15    : DB <=    150    ;
                    16    : DB <=    152    ;
                    17    : DB <=    154    ;
                    18    : DB <=    155    ;
                    19    : DB <=    157    ;
                    20    : DB <=    158    ;
                    21    : DB <=    160    ;
                    22    : DB <=    161    ;
                    23    : DB <=    163    ;
                    24    : DB <=    164    ;
                    25    : DB <=    166    ;
                    26    : DB <=    167    ;
                    27    : DB <=    169    ;
                    28    : DB <=    170    ;
                    29    : DB <=    172    ;
                    30    : DB <=    173    ;
                    31    : DB <=    175    ;
                    32    : DB <=    176    ;
                    33    : DB <=    177    ;
                    34    : DB <=    179    ;
                    35    : DB <=    180    ;
                    36    : DB <=    182    ;
                    37    : DB <=    183    ;
                    38    : DB <=    185    ;
                    39    : DB <=    186    ;
                    40    : DB <=    187    ;
                    41    : DB <=    189    ;
                    42    : DB <=    190    ;
                    43    : DB <=    191    ;
                    44    : DB <=    193    ;
                    45    : DB <=    194    ;
                    46    : DB <=    195    ;
                    47    : DB <=    197    ;
                    48    : DB <=    198    ;
                    49    : DB <=    199    ;
                    50    : DB <=    201    ;
                    51    : DB <=    202    ;
                    52    : DB <=    203    ;
                    53    : DB <=    205    ;
                    54    : DB <=    206    ;
                    55    : DB <=    207    ;
                    56    : DB <=    208    ;
                    57    : DB <=    209    ;
                    58    : DB <=    211    ;
                    59    : DB <=    212    ;
                    60    : DB <=    213    ;
                    61    : DB <=    214    ;
                    62    : DB <=    215    ;
                    63    : DB <=    216    ;
                    64    : DB <=    218    ;
                    65    : DB <=    219    ;
                    66    : DB <=    220    ;
                    67    : DB <=    221    ;
                    68    : DB <=    222    ;
                    69    : DB <=    223    ;
                    70    : DB <=    224    ;
                    71    : DB <=    225    ;
                    72    : DB <=    226    ;
                    73    : DB <=    227    ;
                    74    : DB <=    228    ;
                    75    : DB <=    229    ;
                    76    : DB <=    230    ;
                    77    : DB <=    231    ;
                    78    : DB <=    232    ;
                    79    : DB <=    233    ;
                    80    : DB <=    233    ;
                    81    : DB <=    234    ;
                    82    : DB <=    235    ;
                    83    : DB <=    236    ;
                    84    : DB <=    237    ;
                    85    : DB <=    238    ;
                    86    : DB <=    238    ;
                    87    : DB <=    239    ;
                    88    : DB <=    240    ;
                    89    : DB <=    241    ;
                    90    : DB <=    241    ;
                    91    : DB <=    242    ;
                    92    : DB <=    243    ;
                    93    : DB <=    243    ;
                    94    : DB <=    244    ;
                    95    : DB <=    245    ;
                    96    : DB <=    245    ;
                    97    : DB <=    246    ;
                    98    : DB <=    246    ;
                    99    : DB <=    247    ;
                    100    : DB <=    248    ;
                    101    : DB <=    248    ;
                    102    : DB <=    249    ;
                    103    : DB <=    249    ;
                    104    : DB <=    249    ;
                    105    : DB <=    250    ;
                    106    : DB <=    250    ;
                    107    : DB <=    251    ;
                    108    : DB <=    251    ;
                    109    : DB <=    252    ;
                    110    : DB <=    252    ;
                    111    : DB <=    252    ;
                    112    : DB <=    253    ;
                    113    : DB <=    253    ;
                    114    : DB <=    253    ;
                    115    : DB <=    253    ;
                    116    : DB <=    254    ;
                    117    : DB <=    254    ;
                    118    : DB <=    254    ;
                    119    : DB <=    254    ;
                    120    : DB <=    254    ;
                    121    : DB <=    255    ;
                    122    : DB <=    255    ;
                    123    : DB <=    255    ;
                    124    : DB <=    255    ;
                    125    : DB <=    255    ;
                    126    : DB <=    255    ;
                    127    : DB <=    255    ;
                    128    : DB <=    255    ;
                    129    : DB <=    255    ;
                    130    : DB <=    255    ;
                    131    : DB <=    255    ;
                    132    : DB <=    255    ;
                    133    : DB <=    255    ;
                    134    : DB <=    255    ;
                    135    : DB <=    255    ;
                    136    : DB <=    254    ;
                    137    : DB <=    254    ;
                    138    : DB <=    254    ;
                    139    : DB <=    254    ;
                    140    : DB <=    254    ;
                    141    : DB <=    253    ;
                    142    : DB <=    253    ;
                    143    : DB <=    253    ;
                    144    : DB <=    253    ;
                    145    : DB <=    252    ;
                    146    : DB <=    252    ;
                    147    : DB <=    252    ;
                    148    : DB <=    251    ;
                    149    : DB <=    251    ;
                    150    : DB <=    250    ;
                    151    : DB <=    250    ;
                    152    : DB <=    249    ;
                    153    : DB <=    249    ;
                    154    : DB <=    249    ;
                    155    : DB <=    248    ;
                    156    : DB <=    248    ;
                    157    : DB <=    247    ;
                    158    : DB <=    246    ;
                    159    : DB <=    246    ;
                    160    : DB <=    245    ;
                    161    : DB <=    245    ;
                    162    : DB <=    244    ;
                    163    : DB <=    243    ;
                    164    : DB <=    243    ;
                    165    : DB <=    242    ;
                    166    : DB <=    241    ;
                    167    : DB <=    241    ;
                    168    : DB <=    240    ;
                    169    : DB <=    239    ;
                    170    : DB <=    238    ;
                    171    : DB <=    238    ;
                    172    : DB <=    237    ;
                    173    : DB <=    236    ;
                    174    : DB <=    235    ;
                    175    : DB <=    234    ;
                    176    : DB <=    233    ;
                    177    : DB <=    233    ;
                    178    : DB <=    232    ;
                    179    : DB <=    231    ;
                    180    : DB <=    230    ;
                    181    : DB <=    229    ;
                    182    : DB <=    228    ;
                    183    : DB <=    227    ;
                    184    : DB <=    226    ;
                    185    : DB <=    225    ;
                    186    : DB <=    224    ;
                    187    : DB <=    223    ;
                    188    : DB <=    222    ;
                    189    : DB <=    221    ;
                    190    : DB <=    220    ;
                    191    : DB <=    219    ;
                    192    : DB <=    218    ;
                    193    : DB <=    216    ;
                    194    : DB <=    215    ;
                    195    : DB <=    214    ;
                    196    : DB <=    213    ;
                    197    : DB <=    212    ;
                    198    : DB <=    211    ;
                    199    : DB <=    209    ;
                    200    : DB <=    208    ;
                    201    : DB <=    207    ;
                    202    : DB <=    206    ;
                    203    : DB <=    205    ;
                    204    : DB <=    203    ;
                    205    : DB <=    202    ;
                    206    : DB <=    201    ;
                    207    : DB <=    199    ;
                    208    : DB <=    198    ;
                    209    : DB <=    197    ;
                    210    : DB <=    195    ;
                    211    : DB <=    194    ;
                    212    : DB <=    193    ;
                    213    : DB <=    191    ;
                    214    : DB <=    190    ;
                    215    : DB <=    189    ;
                    216    : DB <=    187    ;
                    217    : DB <=    186    ;
                    218    : DB <=    185    ;
                    219    : DB <=    183    ;
                    220    : DB <=    182    ;
                    221    : DB <=    180    ;
                    222    : DB <=    179    ;
                    223    : DB <=    177    ;
                    224    : DB <=    176    ;
                    225    : DB <=    175    ;
                    226    : DB <=    173    ;
                    227    : DB <=    172    ;
                    228    : DB <=    170    ;
                    229    : DB <=    169    ;
                    230    : DB <=    167    ;
                    231    : DB <=    166    ;
                    232    : DB <=    164    ;
                    233    : DB <=    163    ;
                    234    : DB <=    161    ;
                    235    : DB <=    160    ;
                    236    : DB <=    158    ;
                    237    : DB <=    157    ;
                    238    : DB <=    155    ;
                    239    : DB <=    154    ;
                    240    : DB <=    152    ;
                    241    : DB <=    150    ;
                    242    : DB <=    149    ;
                    243    : DB <=    147    ;
                    244    : DB <=    146    ;
                    245    : DB <=    144    ;
                    246    : DB <=    143    ;
                    247    : DB <=    141    ;
                    248    : DB <=    140    ;
                    249    : DB <=    138    ;
                    250    : DB <=    136    ;
                    251    : DB <=    135    ;
                    252    : DB <=    133    ;
                    253    : DB <=    132    ;
                    254    : DB <=    130    ;
                    255    : DB <=    129    ;
                    256    : DB <=    127    ;
                    257    : DB <=    125    ;
                    258    : DB <=    124    ;
                    259    : DB <=    122    ;
                    260    : DB <=    121    ;
                    261    : DB <=    119    ;
                    262    : DB <=    118    ;
                    263    : DB <=    116    ;
                    264    : DB <=    115    ;
                    265    : DB <=    113    ;
                    266    : DB <=    111    ;
                    267    : DB <=    110    ;
                    268    : DB <=    108    ;
                    269    : DB <=    107    ;
                    270    : DB <=    105    ;
                    271    : DB <=    104    ;
                    272    : DB <=    102    ;
                    273    : DB <=    101    ;
                    274    : DB <=    99    ;
                    275    : DB <=    98    ;
                    276    : DB <=    96    ;
                    277    : DB <=    95    ;
                    278    : DB <=    93    ;
                    279    : DB <=    92    ;
                    280    : DB <=    90    ;
                    281    : DB <=    89    ;
                    282    : DB <=    87    ;
                    283    : DB <=    86    ;
                    284    : DB <=    84    ;
                    285    : DB <=    83    ;
                    286    : DB <=    81    ;
                    287    : DB <=    80    ;
                    288    : DB <=    78    ;
                    289    : DB <=    77    ;
                    290    : DB <=    76    ;
                    291    : DB <=    74    ;
                    292    : DB <=    73    ;
                    293    : DB <=    71    ;
                    294    : DB <=    70    ;
                    295    : DB <=    69    ;
                    296    : DB <=    67    ;
                    297    : DB <=    66    ;
                    298    : DB <=    64    ;
                    299    : DB <=    63    ;
                    300    : DB <=    62    ;
                    301    : DB <=    60    ;
                    302    : DB <=    59    ;
                    303    : DB <=    58    ;
                    304    : DB <=    56    ;
                    305    : DB <=    55    ;
                    306    : DB <=    54    ;
                    307    : DB <=    53    ;
                    308    : DB <=    51    ;
                    309    : DB <=    50    ;
                    310    : DB <=    49    ;
                    311    : DB <=    48    ;
                    312    : DB <=    46    ;
                    313    : DB <=    45    ;
                    314    : DB <=    44    ;
                    315    : DB <=    43    ;
                    316    : DB <=    42    ;
                    317    : DB <=    41    ;
                    318    : DB <=    39    ;
                    319    : DB <=    38    ;
                    320    : DB <=    37    ;
                    321    : DB <=    36    ;
                    322    : DB <=    35    ;
                    323    : DB <=    34    ;
                    324    : DB <=    33    ;
                    325    : DB <=    32    ;
                    326    : DB <=    31    ;
                    327    : DB <=    30    ;
                    328    : DB <=    29    ;
                    329    : DB <=    28    ;
                    330    : DB <=    27    ;
                    331    : DB <=    26    ;
                    332    : DB <=    25    ;
                    333    : DB <=    24    ;
                    334    : DB <=    23    ;
                    335    : DB <=    22    ;
                    336    : DB <=    21    ;
                    337    : DB <=    21    ;
                    338    : DB <=    20    ;
                    339    : DB <=    19    ;
                    340    : DB <=    18    ;
                    341    : DB <=    17    ;
                    342    : DB <=    16    ;
                    343    : DB <=    16    ;
                    344    : DB <=    15    ;
                    345    : DB <=    14    ;
                    346    : DB <=    14    ;
                    347    : DB <=    13    ;
                    348    : DB <=    12    ;
                    349    : DB <=    12    ;
                    350    : DB <=    11    ;
                    351    : DB <=    10    ;
                    352    : DB <=    10    ;
                    353    : DB <=    9    ;
                    354    : DB <=    9    ;
                    355    : DB <=    8    ;
                    356    : DB <=    7    ;
                    357    : DB <=    7    ;
                    358    : DB <=    6    ;
                    359    : DB <=    6    ;
                    360    : DB <=    5    ;
                    361    : DB <=    5    ;
                    362    : DB <=    5    ;
                    363    : DB <=    4    ;
                    364    : DB <=    4    ;
                    365    : DB <=    3    ;
                    366    : DB <=    3    ;
                    367    : DB <=    3    ;
                    368    : DB <=    2    ;
                    369    : DB <=    2    ;
                    370    : DB <=    2    ;
                    371    : DB <=    2    ;
                    372    : DB <=    1    ;
                    373    : DB <=    1    ;
                    374    : DB <=    1    ;
                    375    : DB <=    1    ;
                    376    : DB <=    1    ;
                    377    : DB <=    0    ;
                    378    : DB <=    0    ;
                    379    : DB <=    0    ;
                    380    : DB <=    0    ;
                    381    : DB <=    0    ;
                    382    : DB <=    0    ;
                    383    : DB <=    0    ;
                    384    : DB <=    0    ;
                    385    : DB <=    0    ;
                    386    : DB <=    0    ;
                    387    : DB <=    0    ;
                    388    : DB <=    0    ;
                    389    : DB <=    0    ;
                    390    : DB <=    0    ;
                    391    : DB <=    0    ;
                    392    : DB <=    1    ;
                    393    : DB <=    1    ;
                    394    : DB <=    1    ;
                    395    : DB <=    1    ;
                    396    : DB <=    1    ;
                    397    : DB <=    2    ;
                    398    : DB <=    2    ;
                    399    : DB <=    2    ;
                    400    : DB <=    2    ;
                    401    : DB <=    3    ;
                    402    : DB <=    3    ;
                    403    : DB <=    3    ;
                    404    : DB <=    4    ;
                    405    : DB <=    4    ;
                    406    : DB <=    5    ;
                    407    : DB <=    5    ;
                    408    : DB <=    5    ;
                    409    : DB <=    6    ;
                    410    : DB <=    6    ;
                    411    : DB <=    7    ;
                    412    : DB <=    7    ;
                    413    : DB <=    8    ;
                    414    : DB <=    9    ;
                    415    : DB <=    9    ;
                    416    : DB <=    10    ;
                    417    : DB <=    10    ;
                    418    : DB <=    11    ;
                    419    : DB <=    12    ;
                    420    : DB <=    12    ;
                    421    : DB <=    13    ;
                    422    : DB <=    14    ;
                    423    : DB <=    14    ;
                    424    : DB <=    15    ;
                    425    : DB <=    16    ;
                    426    : DB <=    16    ;
                    427    : DB <=    17    ;
                    428    : DB <=    18    ;
                    429    : DB <=    19    ;
                    430    : DB <=    20    ;
                    431    : DB <=    21    ;
                    432    : DB <=    21    ;
                    433    : DB <=    22    ;
                    434    : DB <=    23    ;
                    435    : DB <=    24    ;
                    436    : DB <=    25    ;
                    437    : DB <=    26    ;
                    438    : DB <=    27    ;
                    439    : DB <=    28    ;
                    440    : DB <=    29    ;
                    441    : DB <=    30    ;
                    442    : DB <=    31    ;
                    443    : DB <=    32    ;
                    444    : DB <=    33    ;
                    445    : DB <=    34    ;
                    446    : DB <=    35    ;
                    447    : DB <=    36    ;
                    448    : DB <=    37    ;
                    449    : DB <=    38    ;
                    450    : DB <=    39    ;
                    451    : DB <=    41    ;
                    452    : DB <=    42    ;
                    453    : DB <=    43    ;
                    454    : DB <=    44    ;
                    455    : DB <=    45    ;
                    456    : DB <=    46    ;
                    457    : DB <=    48    ;
                    458    : DB <=    49    ;
                    459    : DB <=    50    ;
                    460    : DB <=    51    ;
                    461    : DB <=    53    ;
                    462    : DB <=    54    ;
                    463    : DB <=    55    ;
                    464    : DB <=    56    ;
                    465    : DB <=    58    ;
                    466    : DB <=    59    ;
                    467    : DB <=    60    ;
                    468    : DB <=    62    ;
                    469    : DB <=    63    ;
                    470    : DB <=    64    ;
                    471    : DB <=    66    ;
                    472    : DB <=    67    ;
                    473    : DB <=    69    ;
                    474    : DB <=    70    ;
                    475    : DB <=    71    ;
                    476    : DB <=    73    ;
                    477    : DB <=    74    ;
                    478    : DB <=    76    ;
                    479    : DB <=    77    ;
                    480    : DB <=    78    ;
                    481    : DB <=    80    ;
                    482    : DB <=    81    ;
                    483    : DB <=    83    ;
                    484    : DB <=    84    ;
                    485    : DB <=    86    ;
                    486    : DB <=    87    ;
                    487    : DB <=    89    ;
                    488    : DB <=    90    ;
                    489    : DB <=    92    ;
                    490    : DB <=    93    ;
                    491    : DB <=    95    ;
                    492    : DB <=    96    ;
                    493    : DB <=    98    ;
                    494    : DB <=    99    ;
                    495    : DB <=    101    ;
                    496    : DB <=    102    ;
                    497    : DB <=    104    ;
                    498    : DB <=    105    ;
                    499    : DB <=    107    ;
                    500    : DB <=    108    ;
                    501    : DB <=    110    ;
                    502    : DB <=    111    ;
                    503    : DB <=    113    ;
                    504    : DB <=    115    ;
                    505    : DB <=    116    ;
                    506    : DB <=    118    ;
                    507    : DB <=    119    ;
                    508    : DB <=    121    ;
                    509    : DB <=    122    ;
                    510    : DB <=    124    ;
                    511    : DB <=    125    ;
                endcase
                horizontalCount <= horizontalCount + 1;
                end
                
            // square        
            2'b01:
                begin
                    if ( DB >= 1 && DB <= 254 ) begin
                        DB <= 0;
                    end
                    if ( horizontalCount % 256 == 0 ) begin
                        DB <= 255 - DB;
                    end
                    horizontalCount <= horizontalCount + 1;
                end
           
           // triangle
            2'b10: 
                begin 
                    if ( DB == 255 - 1  ) begin
                        upDownFlag <= 1;
                    end
                    else if ( DB == 0 + 1 ) begin 
                        upDownFlag <= 0;
                    end
                    if ( upDownFlag == 0 ) begin
                        DB <= DB + 1;
                    end
                    else if ( upDownFlag == 1 ) begin
                        DB <= DB - 1;
                    end
                end     
                              
            2'b11: // sawtooth
                begin
                    DB <= DB + 1;
                end        
        endcase
        end
    end
    
endmodule
